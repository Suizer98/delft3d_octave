// For discussion on this netCDF format please refer to:
// http://public.deltares.nl/display/NETCDF/netCDF
netCDF runid_his.nc {
dimensions:
	time = UNLIMITED ; (3601 currently)
	stations = 6 ;
	station_name_len = 40 ;

variables:
	// Preference 'PRESERVE_FVD':  false,
	// dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
	double station_x_coordinate(stations), shape = [6]
		station_x_coordinate:units = "m" ;
		station_x_coordinate:standard_name = "projection_x_coordinate" ;
		station_x_coordinate:long_name = "x" ;
	double station_y_coordinate(stations), shape = [6]
		station_y_coordinate:units = "m" ;
		station_y_coordinate:standard_name = "projection_y_coordinate" ;
		station_y_coordinate:long_name = "y" ;
	char station_id(stations,station_name_len), shape = [6 40]
		station_id:cf_role = "timeseries_id" ;
		station_id:long_name = "Observation station identifier" ;
	char station_name(stations,station_name_len), shape = [6 40]
		station_name:cf_role = "timeseries_id" ;
		station_name:long_name = "Observation station name" ;
	double waterlevel(time,stations), shape = [3601 6]
		waterlevel:standard_name = "sea_surface_height" ;
		waterlevel:long_name = "Water level" ;
		waterlevel:units = "m" ;
		waterlevel:coordinates = "station_x_coordinate station_y_coordinate station_name" ;
		waterlevel:_FillValue = -999 ;
	double x_velocity(time,stations), shape = [3601 6]
		x_velocity:standard_name = "eastward_sea_water_velocity" ;
		x_velocity:long_name = "Horizontal/eastward component of cell center velocity vector." ;
		x_velocity:units = "m s-1" ;
		x_velocity:coordinates = "station_x_coordinate station_y_coordinate station_name" ;
		x_velocity:_FillValue = -999 ;
	double y_velocity(time,stations), shape = [3601 6]
		y_velocity:standard_name = "northward_sea_water_velocity" ;
		y_velocity:long_name = "Vertical/northward component of cell center velocity vector." ;
		y_velocity:units = "m s-1" ;
		y_velocity:coordinates = "station_x_coordinate station_y_coordinate station_name" ;
		y_velocity:_FillValue = -999 ;
	double time(time), shape = [3601]
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;

//global attributes:
		:institution = "Deltares" ;
		:references = "http://www.deltares.nl" ;
		:source = "Deltares, D-Flow FM Version 1.1.72.000000, Jul 11 2013, 20:09:35, model" ;
		:history = "Created on 2013-07-18T23:22:39+0200, D-Flow FM" ;
		:Conventions = "CF-1.5:Deltares-0.1" ;

}
