// The netCDF-CF conventions for grids are defined here:
// http://cf-pcmdi.llnl.gov/documents/cf-conventions/
// This grid file can be loaded into matlab with QuickPlot (d3d_qp.m) and ADAGUC.knmi.nl.
// To create this netCDF file with Matlab please see ncwritetutorial_grid_lat_lon_swath
NetCDF-3 Classic ncwritetutorial_grid_lat_lon_swath.nc {

  dimensions:
    NUMCELLS = 3 ;
    NUMROWS = 5 ;
    bounds = 4 ;

  variables:
    // Preference 'PRESERVE_FVD':  false,
    // dimensions consistent with ncBrowse, not with native MATLAB netcdf package.
    double time(NUMROWS,NUMCELLS), shape = [5 3]
      :standard_name = "time" 
      :long_name = "time" 
      :units = "days since 1970-01-01 00:00:00+08:00" 
      :axis = "T" 
    double lon(NUMROWS,NUMCELLS), shape = [5 3]
      :standard_name = "longitude" 
      :long_name = "Longitude" 
      :units = "degrees_east" 
      :axis = "X" 
      :_FillValue = NaN 
      :grid_mapping = "wgs84" 
      :actual_range = 2 6 
      :bounds = "lon_bnds" 
    double lat(NUMROWS,NUMCELLS), shape = [5 3]
      :standard_name = "latitude" 
      :long_name = "Latitude" 
      :units = "degrees_north" 
      :axis = "Y" 
      :_FillValue = NaN 
      :grid_mapping = "wgs84" 
      :actual_range = 50 54 
      :bounds = "lat_bnds" 
    int32 wgs84([]), shape = [1]
      :name = "WGS 84" 
      :epsg = 4326 
      :grid_mapping_name = "latitude_longitude" 
      :semi_major_axis = 6.37814e+06 
      :semi_minor_axis = 6.35675e+06 
      :inverse_flattening = 298.257 
      :comment = "value is equal to EPSG code" 
      :proj4_params = "+proj=longlat +ellps=WGS84 +datum=WGS84 +no_defs" 
      :projection_name = "Latitude Longitude" 
      :EPSG_code = "EPSG:4326" 
    double lon_bnds(NUMROWS,NUMCELLS,bounds), shape = [5 3 4]
      :standard_name = "longitude" 
      :long_name = "Longitude bounds" 
      :units = "degrees_east" 
      :_FillValue = NaN 
      :actual_range = 1 7 
    double lat_bnds(NUMROWS,NUMCELLS,bounds), shape = [5 3 4]
      :standard_name = "latitude" 
      :long_name = "Latitude bounds" 
      :units = "degrees_north" 
      :_FillValue = NaN 
      :actual_range = 49.5 54.5 
    double depth(NUMROWS,NUMCELLS), shape = [5 3]
      :standard_name = "sea_floor_depth_below_geoid" 
      :long_name = "bottom depth" 
      :units = "m" 
      :_FillValue = NaN 
      :actual_range = 1 114 
      :grid_mapping = "wgs84" 
      :coordinates = "lat lon" 

  //global Attributes:
      :title = "ncwritetutorial_grid_lat_lon_swath" 
      :institution = "Deltares" 
      :source = "" 
      :history = "$HeadURL: https://svn.oss.deltares.nl/repos/openearthtools/trunk/matlab/io/netcdf/nctools/ncwritetutorial_grid_lat_lon_curvilinear.m $ $Id: ncwritetutorial_grid_lat_lon_curvilinear.m 8831 2013-06-19 08:05:18Z boer_g $" 
      :references = "http://svn.oss.deltares.nl" 
      :email = "" 
      :featureType = "grid" 
      :comment = "" 
      :version = "" 
      :Conventions = "CF-1.6" 
      :terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: Deltares" 
      :disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." 
      :time_coverage_start = "2000-01-01T00:00" 
      :time_coverage_end = "2000-01-01T00:00" 


}
