netcdf dgC_his {
dimensions:
	time = 1003 ;
	Layer = 40 ;
	LayerInterf = 41 ;
	Fraction = 1 ;
	bounds2 = 2 ;
	platform_name_len = 20 ;
	Station = 152 ;
	crs_name_len = 20 ;
	Crosssection = 18 ;
	start_end = 2 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1970-01-01 00:00:00 " ;
		time:axis = "T" ;
		time:actual_range = "2002-05-26 10:00:00\t2002-06-02 09:00:00" ;
	char platform_name(Station, platform_name_len) ;
		platform_name:standard_name = "platform_name" ;
		platform_name:long_name = "Name of monitoring station" ;
		platform_name:delft3d_name = "NAMST" ;
		platform_name:cf_role = "timeseries_id" ;
	float platform_m_index(Station) ;
		platform_m_index:long_name = "Delft3D-FLOW m index of station" ;
		platform_m_index:units = "1" ;
		platform_m_index:delft3d_name = "MNSTAT" ;
		platform_m_index:_FillValue = -1.#IND00f ;
		platform_m_index:actual_range = 3., 138. ;
	float platform_n_index(Station) ;
		platform_n_index:long_name = "Delft3D-FLOW n index of station" ;
		platform_n_index:units = "1" ;
		platform_n_index:delft3d_name = "MNSTAT" ;
		platform_n_index:_FillValue = -1.#IND00f ;
		platform_n_index:actual_range = 7., 34. ;
	float platform_angle(Station) ;
		platform_angle:long_name = "Orientation ksi-axis w.r.t. pos.x-axis at water level point" ;
		platform_angle:delft3d_name = "ALFAS" ;
	char crs_name(Crosssection, crs_name_len) ;
		crs_name:standard_name = "platform_name" ;
		crs_name:long_name = "Name of monitoring cross-section" ;
		crs_name:delft3d_name = "NAMTRA" ;
		crs_name:cf_role = "timeseries_id" ;
	float crs_m(Crosssection, start_end) ;
		crs_m:long_name = "Delft3D-FLOW m indices of cross-section" ;
		crs_m:units = "1" ;
		crs_m:delft3d_name = "MNTRA" ;
		crs_m:_FillValue = -1.#IND00f ;
		crs_m:actual_range = 9., 138. ;
	float crs_n(Crosssection, start_end) ;
		crs_n:long_name = "Delft3D-FLOW n indices of cross-section" ;
		crs_n:units = "1" ;
		crs_n:delft3d_name = "MNTRA" ;
		crs_n:_FillValue = -1.#IND00f ;
		crs_n:actual_range = 3., 33. ;
	float x(Station) ;
		x:standard_name = "projection_x_coordinate" ;
		x:long_name = "x of station" ;
		x:units = "m" ;
		x:axis = "X" ;
		x:delft3d_name = "XYSTAT" ;
		x:_FillValue = -1.#IND00f ;
		x:actual_range = 75745.53125, 77579.96875 ;
	float y(Station) ;
		y:standard_name = "projection_y_coordinate" ;
		y:long_name = "y of station" ;
		y:units = "m" ;
		y:axis = "Y" ;
		y:delft3d_name = "XYSTAT" ;
		y:_FillValue = -1.#IND00f ;
		y:actual_range = 366566.40625, 369509.53125 ;
	float longitude(Station) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "Longitude of station" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:delft3d_name = "XYSTAT" ;
		longitude:_FillValue = -1.#IND00f ;
		longitude:actual_range = 4.25119459783757, 4.27686155660913 ;
	float latitude(Station) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "Latitude of station" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:delft3d_name = "XYSTAT" ;
		latitude:_FillValue = -1.#IND00f ;
		latitude:actual_range = 51.2828413546755, 51.30947637028 ;
	float crs_x(Crosssection) ;
		crs_x:standard_name = "projection_x_coordinate" ;
		crs_x:long_name = "x of cross-section" ;
		crs_x:units = "m" ;
		crs_x:axis = "X" ;
		crs_x:delft3d_name = "XYTRA" ;
		crs_x:_FillValue = -1.#IND00f ;
		crs_x:actual_range = 75602.375, 77217.2734375 ;
	float crs_y(Crosssection) ;
		crs_y:standard_name = "projection_y_coordinate" ;
		crs_y:long_name = "y of cross-section" ;
		crs_y:units = "m" ;
		crs_y:axis = "Y" ;
		crs_y:delft3d_name = "XYTRA" ;
		crs_y:_FillValue = -1.#IND00f ;
		crs_y:actual_range = 366566.40625, 369509.53125 ;
	float crs_longitude(Crosssection, start_end) ;
		crs_longitude:standard_name = "longitude" ;
		crs_longitude:long_name = "Longitude of cross-section" ;
		crs_longitude:units = "degrees_east" ;
		crs_longitude:axis = "X" ;
		crs_longitude:delft3d_name = "XYTRA" ;
		crs_longitude:_FillValue = -1.#IND00f ;
		crs_longitude:actual_range = 4.24912241693128, 4.27189634614567 ;
	float crs_latitude(Crosssection, start_end) ;
		crs_latitude:standard_name = "latitude" ;
		crs_latitude:long_name = "Latitude of cross-section" ;
		crs_latitude:units = "degrees_north" ;
		crs_latitude:axis = "Y" ;
		crs_latitude:delft3d_name = "XYTRA" ;
		crs_latitude:_FillValue = -1.#IND00f ;
		crs_latitude:actual_range = 51.2817788284517, 51.3085817491024 ;
	float Layer(Layer) ;
		Layer:long_name = "sigma at layer midpoints" ;
		Layer:standard_name = "ocean_sigma_coordinate" ;
		Layer:positive = "up" ;
		Layer:actual_range = -0.999666506308131, -0.0632033199071884 ;
		Layer:formula_terms = "sigma: Layer eta: waterlevel depth: depth" ;
		Layer:comment = "The surface layer has index k=1 and is sigma=0, the bottom layer has index kmax and is sigma=-1." ;
		Layer:delft3d_name = "his-const:KMAX his-const:LAYER_MODEL his-const:THICK" ;
	float LayerInterf(LayerInterf) ;
		LayerInterf:long_name = "sigma at layer interfaces" ;
		LayerInterf:standard_name = "ocean_sigma_coordinate" ;
		LayerInterf:positive = "up" ;
		LayerInterf:actual_range = -1.00000001327135, 0. ;
		LayerInterf:formula_terms = "sigma: LayerInterf eta: waterlevel depth: depth" ;
		LayerInterf:comment = "The surface layer has index k=1 and is sigma=0, the bottom layer has index kmax and is sigma=-1." ;
		LayerInterf:delft3d_name = "his-const:KMAX his-const:LAYER_MODEL his-const:THICK" ;
	float depth(Station) ;
		depth:standard_name = "altitude" ;
		depth:long_name = "Depth in station" ;
		depth:units = "m" ;
		depth:positive = "down" ;
		depth:coordinates = "x y platform_name" ;
		depth:delft3d_name = "DPS" ;
		depth:comment = "" ;
		depth:actual_range = 0.162000000476837, 16.942455291748 ;
	float waterlevel(time, Station) ;
		waterlevel:standard_name = "sea_surface_elevation" ;
		waterlevel:long_name = "Water-level in station (zeta point)" ;
		waterlevel:units = "m" ;
		waterlevel:positive = "up" ;
		waterlevel:coordinates = "x y platform_name" ;
		waterlevel:delft3d_name = "ZWL" ;
		waterlevel:_FillValue = -1.#IND00f ;
		waterlevel:actual_range = -0.460175931453705, 5.84168863296509 ;
	single mask(time,Station), shape = [3803 150]
		mask:standard_name = "" ;
		mask:long_name = "active" ;
		mask:units = "1" ;
		mask:coordinates = "latitude longitude platform_name" ;
		mask:delft3d_name = "ZKFS" ;
		mask:_FillValue = NaN f;
		mask:actual_range = 0 1 ;
		mask:flag_values = 0 1 ;
		mask:flag_meanings = "inactive active " ;
	float u_x(time, Station, Layer) ;
		u_x:standard_name = "sea_water_x_velocity" ;
		u_x:long_name = "velocity, x-component" ;
		u_x:units = "m/s" ;
		u_x:coordinates = "x y platform_name" ;
		u_x:delft3d_name = "ZCURU" ;
		u_x:_FillValue = -1.#IND00f ;
		u_x:actual_range = -0.973308503627777, 1.31783068180084 ;
	float u_y(time, Station, Layer) ;
		u_y:standard_name = "sea_water_y_velocity" ;
		u_y:long_name = "velocity, y-component" ;
		u_y:units = "m/s" ;
		u_y:coordinates = "x y platform_name" ;
		u_y:delft3d_name = "ZCURV" ;
		u_y:_FillValue = -1.#IND00f ;
		u_y:actual_range = -0.92728465795517, 0.715223848819733 ;
	float u_z(time, Station, Layer) ;
		u_z:standard_name = "upward_sea_water_velocity" ;
		u_z:long_name = "velocity, z-component" ;
		u_z:units = "m/s" ;
		u_z:positive = "up" ;
		u_z:coordinates = "x y platform_name" ;
		u_z:delft3d_name = "ZCURW" ;
		u_z:_FillValue = -1.#IND00f ;
		u_z:actual_range = -0.177295297384262, 0.257271468639374 ;
	float Q(time, Crosssection) ;
		Q:standard_name = "water_flux_into_sea_water" ;
		Q:long_name = "Monumentary discharge through cross section (velocity points)" ;
		Q:units = "m3/s" ;
		Q:coordinates = "crs_x crs_y crs_name" ;
		Q:delft3d_name = "CTR" ;
		Q:_FillValue = -1.#IND00f ;
		Q:actual_range = 1.#INF0000000000, -1.#INF0000000000 ;
	float CQ(time, Crosssection) ;
		CQ:standard_name = "water_flux_into_sea_water" ;
		CQ:long_name = "Total discharge through cross section (velocity points)" ;
		CQ:units = "m3" ;
		CQ:coordinates = "crs_x crs_y crs_name" ;
		CQ:delft3d_name = "FLTR" ;
		CQ:_FillValue = -1.#IND00f ;
		CQ:actual_range = -72419024., 13368214. ;
	float tau_x(time, Station) ;
		tau_x:standard_name = "surface_downward_x_stress" ;
		tau_x:long_name = "Bottom stress U in station (zeta point)" ;
		tau_x:units = "N m-2" ;
		tau_x:coordinates = "x y platform_name" ;
		tau_x:delft3d_name = "ZTAUKS" ;
		tau_x:_FillValue = -1.#IND00f ;
		tau_x:actual_range = -2.35219240188599, 3.14754724502563 ;
		tau_x:comment = "The bed shear stresses are in real world directions x and y" ;
	float tau_y(time, Station) ;
		tau_y:standard_name = "surface_downward_y_stress" ;
		tau_y:long_name = "Bottom stress V in station (zeta point)" ;
		tau_y:units = "N m-2" ;
		tau_y:coordinates = "x y platform_name" ;
		tau_y:delft3d_name = "ZTAUET" ;
		tau_y:_FillValue = -1.#IND00f ;
		tau_y:actual_range = -1.23002445697784, 2.36216640472412 ;
		tau_y:comment = "The bed shear stresses are in real world directions x and y" ;
	float density(time, Station, Layer) ;
		density:standard_name = "sea_water_density" ;
		density:long_name = "Density in station" ;
		density:units = "kg/m3" ;
		density:coordinates = "x y platform_name" ;
		density:delft3d_name = "ZRHO" ;
		density:_FillValue = -1.#IND00f ;
		density:actual_range = 1004.97137451172, 1008.29388427734 ;
	float salinity(time, Station, Layer) ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:long_name = "Salinity in station" ;
		salinity:units = "psu" ;
		salinity:coordinates = "x y platform_name" ;
		salinity:delft3d_name = "GRO" ;
		salinity:_FillValue = -1.#IND00f ;
		salinity:actual_range = 7.75254106521606, 11.8001956939697 ;
	single temperature(time,Station,Layer), shape = [3803 150 10]
		temperature:standard_name = "sea_water_temperature" ;
		temperature:long_name = "Temperature in station" ;
		temperature:units = "degree_Celsius" ;
		temperature:coordinates = "latitude longitude platform_name" ;
		temperature:delft3d_name = "GRO" ;
		temperature:_FillValue = NaN f;
		temperature:actual_range = -0.00931975 11.8603 ;
	float sediment_coh(time, Station, Layer) ;
		sediment_coh:standard_name = "concentration_of_suspended_matter_in_sea_water" ;
		sediment_coh:long_name = "Concentration of sediment_coh per layer in station" ;
		sediment_coh:units = "kg/m3" ;
		sediment_coh:coordinates = "x y platform_name" ;
		sediment_coh:delft3d_name = "GRO" ;
		sediment_coh:_FillValue = -1.#IND00f ;
		sediment_coh:actual_range = -0.00832465570420027, 2.26311326026917 ;
	float tke(time, Station, LayerInterf) ;
		tke:standard_name = "specific_kinetic_energy_of_sea_water" ;
		tke:long_name = "Turbulent kinetic energy in station" ;
		tke:units = "m2/s2" ;
		tke:coordinates = "x y platform_name" ;
		tke:delft3d_name = "ZTUR" ;
		tke:_FillValue = -1.#IND00f ;
		tke:actual_range = 0., 0.0482837557792664 ;
	float eps(time, Station, LayerInterf) ;
		eps:standard_name = "ocean_kinetic_energy_dissipation_per_unit_area_due_to_vertical_friction" ;
		eps:long_name = "Turbulent dissipation in station" ;
		eps:units = "m2/s3" ;
		eps:coordinates = "x y platform_name" ;
		eps:delft3d_name = "ZTUR" ;
		eps:_FillValue = -1.#IND00f ;
		eps:actual_range = 0., 0.798907995223999 ;
	float viscosity_z(time, Station, LayerInterf) ;
		viscosity_z:standard_name = "ocean_vertical_momentum_diffusivity" ;
		viscosity_z:long_name = "Vertical eddy viscosity-3D" ;
		viscosity_z:units = "m^2/s" ;
		viscosity_z:coordinates = "x y platform_name" ;
		viscosity_z:delft3d_name = "ZVICWW" ;
		viscosity_z:_FillValue = -1.#IND00f ;
		viscosity_z:actual_range = 0., 0.169904321432114 ;
	float diffusivity_z(time, Station, LayerInterf) ;
		diffusivity_z:standard_name = "ocean_vertical_tracer_diffusivity" ;
		diffusivity_z:long_name = "Vertical eddy diffusivity-3D" ;
		diffusivity_z:units = "m^2/s" ;
		diffusivity_z:coordinates = "x y platform_name" ;
		diffusivity_z:delft3d_name = "ZDICWW" ;
		diffusivity_z:_FillValue = -1.#IND00f ;
		diffusivity_z:actual_range = 0., 0.169904321432114 ;
	float Ri(time, Station, LayerInterf) ;
		Ri:standard_name = "richardson_number_in_sea_water" ;
		Ri:long_name = "Richardson number" ;
		Ri:units = "-" ;
		Ri:coordinates = "x y platform_name" ;
		Ri:delft3d_name = "ZRICH" ;
		Ri:_FillValue = -1.#IND00f ;
		Ri:actual_range = -42776.19921875, 141448.875 ;
	float morphological_depth(time, Station) ;
		morphological_depth:standard_name = "" ;
		morphological_depth:long_name = "Morphological depth at station (zeta point)" ;
		morphological_depth:units = "m" ;
		morphological_depth:coordinates = "x y platform_name" ;
		morphological_depth:delft3d_name = "ZDPS" ;
		morphological_depth:_FillValue = -1.#IND00f ;
		morphological_depth:actual_range = 0.155364751815796, 16.9475440979004 ;
	float available_mass_of_sediment(time, Station, Fraction) ;
		available_mass_of_sediment:standard_name = "" ;
		available_mass_of_sediment:long_name = "Available mass of sediment at bed at station" ;
		available_mass_of_sediment:units = "kg/m2" ;
		available_mass_of_sediment:coordinates = "x y platform_name" ;
		available_mass_of_sediment:delft3d_name = "ZBDSED" ;
		available_mass_of_sediment:_FillValue = -1.#IND00f ;
		available_mass_of_sediment:actual_range = -4.13602379012445e-007, 58.5657653808594 ;
	float bed_load_transport(time, Crosssection, Fraction) ;
		bed_load_transport:standard_name = "" ;
		bed_load_transport:long_name = "Momentary bed load transport through section" ;
		bed_load_transport:units = "m3/s" ;
		bed_load_transport:coordinates = "crs_x crs_y crs_name" ;
		bed_load_transport:delft3d_name = "SBTR" ;
		bed_load_transport:_FillValue = -1.#IND00f ;
		bed_load_transport:actual_range = 0., 0. ;
	float cumulative_bed_load_transport(time, Crosssection, Fraction) ;
		cumulative_bed_load_transport:standard_name = "" ;
		cumulative_bed_load_transport:long_name = "Cumulative bed load transport through section" ;
		cumulative_bed_load_transport:units = "m3" ;
		cumulative_bed_load_transport:coordinates = "crs_x crs_y crs_name" ;
		cumulative_bed_load_transport:delft3d_name = "SBTRC" ;
		cumulative_bed_load_transport:_FillValue = -1.#IND00f ;
		cumulative_bed_load_transport:actual_range = 0., 0. ;
	float suspended_load_transport(time, Crosssection, Fraction) ;
		suspended_load_transport:standard_name = "" ;
		suspended_load_transport:long_name = "Momentary susp. load transport through section" ;
		suspended_load_transport:units = "m3/s" ;
		suspended_load_transport:coordinates = "crs_x crs_y crs_name" ;
		suspended_load_transport:delft3d_name = "SSTR" ;
		suspended_load_transport:_FillValue = -1.#IND00f ;
		suspended_load_transport:actual_range = -0.0500059761106968, 0.143801242113113 ;
	float cumulative_suspended_load_transport(time, Crosssection, Fraction) ;
		cumulative_suspended_load_transport:standard_name = "" ;
		cumulative_suspended_load_transport:long_name = "Cumulative susp. load transport through section" ;
		cumulative_suspended_load_transport:units = "m3" ;
		cumulative_suspended_load_transport:coordinates = "crs_x crs_y crs_name" ;
		cumulative_suspended_load_transport:delft3d_name = "SSTRC" ;
		cumulative_suspended_load_transport:_FillValue = -1.#IND00f ;
		cumulative_suspended_load_transport:actual_range = -1005.068359375, 3350.57495117188 ;

// global attributes:
		:title = "" ;
		:institution = "" ;
		:source = "Delft3D trih file" ;
		:history = "Original filename: trih-RUNID.dat, Deltares, FLOW2D3D Version X, DATE, file version: X, file date: DATA, transformation to netCDF: HeadURL Id" ;
		:references = "http://svn.oss.deltares.nl" ;
		:email = "" ;
		:comment = "" ;
		:version = "" ;
		:Conventions = "CF-1.6" ;
		:terms_for_use = "These data can be used freely for research purposes provided that the following source is acknowledged: " ;
		:disclaimer = "This data is made available in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE." ;
		:delft3d_description = "                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"                              \n",
			"" ;
		:time_coverage_start = "yyyy-mm-ddTHH:00" ;
		:time_coverage_end = "yyyy-mm-ddTHH:00" ;
		:featureType = "timeSeries" ;
}
